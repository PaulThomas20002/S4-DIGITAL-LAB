module not_gate(x,z);
  input x;
  output z;
  not gl(z,x);
endmodule
